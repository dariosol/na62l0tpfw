  --Example instantiation for system 'nios'
  nios_inst : nios
    port map(
      s_address_from_the_iobusMAC_0 => s_address_from_the_iobusMAC_0,
      s_address_from_the_iobusMAC_1 => s_address_from_the_iobusMAC_1,
      s_address_from_the_iobusMAC_2 => s_address_from_the_iobusMAC_2,
      s_address_from_the_iobusMAC_3 => s_address_from_the_iobusMAC_3,
      s_address_from_the_iobusMAC_4 => s_address_from_the_iobusMAC_4,
      s_address_from_the_iobusMAC_5 => s_address_from_the_iobusMAC_5,
      s_address_from_the_iobusMAC_6 => s_address_from_the_iobusMAC_6,
      s_address_from_the_iobusMAC_7 => s_address_from_the_iobusMAC_7,
      s_address_from_the_iobusMDIO_0 => s_address_from_the_iobusMDIO_0,
      s_address_from_the_iobusMDIO_1 => s_address_from_the_iobusMDIO_1,
      s_address_from_the_iobusMDIO_2 => s_address_from_the_iobusMDIO_2,
      s_address_from_the_iobusMDIO_3 => s_address_from_the_iobusMDIO_3,
      s_address_from_the_iobusMDIO_4 => s_address_from_the_iobusMDIO_4,
      s_address_from_the_iobusMDIO_5 => s_address_from_the_iobusMDIO_5,
      s_address_from_the_iobusMDIO_6 => s_address_from_the_iobusMDIO_6,
      s_address_from_the_iobusMDIO_7 => s_address_from_the_iobusMDIO_7,
      s_address_from_the_iobusREGFILE_0 => s_address_from_the_iobusREGFILE_0,
      s_clk_from_the_iobusMAC_0 => s_clk_from_the_iobusMAC_0,
      s_clk_from_the_iobusMAC_1 => s_clk_from_the_iobusMAC_1,
      s_clk_from_the_iobusMAC_2 => s_clk_from_the_iobusMAC_2,
      s_clk_from_the_iobusMAC_3 => s_clk_from_the_iobusMAC_3,
      s_clk_from_the_iobusMAC_4 => s_clk_from_the_iobusMAC_4,
      s_clk_from_the_iobusMAC_5 => s_clk_from_the_iobusMAC_5,
      s_clk_from_the_iobusMAC_6 => s_clk_from_the_iobusMAC_6,
      s_clk_from_the_iobusMAC_7 => s_clk_from_the_iobusMAC_7,
      s_clk_from_the_iobusMDIO_0 => s_clk_from_the_iobusMDIO_0,
      s_clk_from_the_iobusMDIO_1 => s_clk_from_the_iobusMDIO_1,
      s_clk_from_the_iobusMDIO_2 => s_clk_from_the_iobusMDIO_2,
      s_clk_from_the_iobusMDIO_3 => s_clk_from_the_iobusMDIO_3,
      s_clk_from_the_iobusMDIO_4 => s_clk_from_the_iobusMDIO_4,
      s_clk_from_the_iobusMDIO_5 => s_clk_from_the_iobusMDIO_5,
      s_clk_from_the_iobusMDIO_6 => s_clk_from_the_iobusMDIO_6,
      s_clk_from_the_iobusMDIO_7 => s_clk_from_the_iobusMDIO_7,
      s_clk_from_the_iobusREGFILE_0 => s_clk_from_the_iobusREGFILE_0,
      s_read_from_the_iobusMAC_0 => s_read_from_the_iobusMAC_0,
      s_read_from_the_iobusMAC_1 => s_read_from_the_iobusMAC_1,
      s_read_from_the_iobusMAC_2 => s_read_from_the_iobusMAC_2,
      s_read_from_the_iobusMAC_3 => s_read_from_the_iobusMAC_3,
      s_read_from_the_iobusMAC_4 => s_read_from_the_iobusMAC_4,
      s_read_from_the_iobusMAC_5 => s_read_from_the_iobusMAC_5,
      s_read_from_the_iobusMAC_6 => s_read_from_the_iobusMAC_6,
      s_read_from_the_iobusMAC_7 => s_read_from_the_iobusMAC_7,
      s_read_from_the_iobusMDIO_0 => s_read_from_the_iobusMDIO_0,
      s_read_from_the_iobusMDIO_1 => s_read_from_the_iobusMDIO_1,
      s_read_from_the_iobusMDIO_2 => s_read_from_the_iobusMDIO_2,
      s_read_from_the_iobusMDIO_3 => s_read_from_the_iobusMDIO_3,
      s_read_from_the_iobusMDIO_4 => s_read_from_the_iobusMDIO_4,
      s_read_from_the_iobusMDIO_5 => s_read_from_the_iobusMDIO_5,
      s_read_from_the_iobusMDIO_6 => s_read_from_the_iobusMDIO_6,
      s_read_from_the_iobusMDIO_7 => s_read_from_the_iobusMDIO_7,
      s_read_from_the_iobusREGFILE_0 => s_read_from_the_iobusREGFILE_0,
      s_rst_from_the_iobusMAC_0 => s_rst_from_the_iobusMAC_0,
      s_rst_from_the_iobusMAC_1 => s_rst_from_the_iobusMAC_1,
      s_rst_from_the_iobusMAC_2 => s_rst_from_the_iobusMAC_2,
      s_rst_from_the_iobusMAC_3 => s_rst_from_the_iobusMAC_3,
      s_rst_from_the_iobusMAC_4 => s_rst_from_the_iobusMAC_4,
      s_rst_from_the_iobusMAC_5 => s_rst_from_the_iobusMAC_5,
      s_rst_from_the_iobusMAC_6 => s_rst_from_the_iobusMAC_6,
      s_rst_from_the_iobusMAC_7 => s_rst_from_the_iobusMAC_7,
      s_rst_from_the_iobusMDIO_0 => s_rst_from_the_iobusMDIO_0,
      s_rst_from_the_iobusMDIO_1 => s_rst_from_the_iobusMDIO_1,
      s_rst_from_the_iobusMDIO_2 => s_rst_from_the_iobusMDIO_2,
      s_rst_from_the_iobusMDIO_3 => s_rst_from_the_iobusMDIO_3,
      s_rst_from_the_iobusMDIO_4 => s_rst_from_the_iobusMDIO_4,
      s_rst_from_the_iobusMDIO_5 => s_rst_from_the_iobusMDIO_5,
      s_rst_from_the_iobusMDIO_6 => s_rst_from_the_iobusMDIO_6,
      s_rst_from_the_iobusMDIO_7 => s_rst_from_the_iobusMDIO_7,
      s_rst_from_the_iobusREGFILE_0 => s_rst_from_the_iobusREGFILE_0,
      s_write_from_the_iobusMAC_0 => s_write_from_the_iobusMAC_0,
      s_write_from_the_iobusMAC_1 => s_write_from_the_iobusMAC_1,
      s_write_from_the_iobusMAC_2 => s_write_from_the_iobusMAC_2,
      s_write_from_the_iobusMAC_3 => s_write_from_the_iobusMAC_3,
      s_write_from_the_iobusMAC_4 => s_write_from_the_iobusMAC_4,
      s_write_from_the_iobusMAC_5 => s_write_from_the_iobusMAC_5,
      s_write_from_the_iobusMAC_6 => s_write_from_the_iobusMAC_6,
      s_write_from_the_iobusMAC_7 => s_write_from_the_iobusMAC_7,
      s_write_from_the_iobusMDIO_0 => s_write_from_the_iobusMDIO_0,
      s_write_from_the_iobusMDIO_1 => s_write_from_the_iobusMDIO_1,
      s_write_from_the_iobusMDIO_2 => s_write_from_the_iobusMDIO_2,
      s_write_from_the_iobusMDIO_3 => s_write_from_the_iobusMDIO_3,
      s_write_from_the_iobusMDIO_4 => s_write_from_the_iobusMDIO_4,
      s_write_from_the_iobusMDIO_5 => s_write_from_the_iobusMDIO_5,
      s_write_from_the_iobusMDIO_6 => s_write_from_the_iobusMDIO_6,
      s_write_from_the_iobusMDIO_7 => s_write_from_the_iobusMDIO_7,
      s_write_from_the_iobusREGFILE_0 => s_write_from_the_iobusREGFILE_0,
      s_writedata_from_the_iobusMAC_0 => s_writedata_from_the_iobusMAC_0,
      s_writedata_from_the_iobusMAC_1 => s_writedata_from_the_iobusMAC_1,
      s_writedata_from_the_iobusMAC_2 => s_writedata_from_the_iobusMAC_2,
      s_writedata_from_the_iobusMAC_3 => s_writedata_from_the_iobusMAC_3,
      s_writedata_from_the_iobusMAC_4 => s_writedata_from_the_iobusMAC_4,
      s_writedata_from_the_iobusMAC_5 => s_writedata_from_the_iobusMAC_5,
      s_writedata_from_the_iobusMAC_6 => s_writedata_from_the_iobusMAC_6,
      s_writedata_from_the_iobusMAC_7 => s_writedata_from_the_iobusMAC_7,
      s_writedata_from_the_iobusMDIO_0 => s_writedata_from_the_iobusMDIO_0,
      s_writedata_from_the_iobusMDIO_1 => s_writedata_from_the_iobusMDIO_1,
      s_writedata_from_the_iobusMDIO_2 => s_writedata_from_the_iobusMDIO_2,
      s_writedata_from_the_iobusMDIO_3 => s_writedata_from_the_iobusMDIO_3,
      s_writedata_from_the_iobusMDIO_4 => s_writedata_from_the_iobusMDIO_4,
      s_writedata_from_the_iobusMDIO_5 => s_writedata_from_the_iobusMDIO_5,
      s_writedata_from_the_iobusMDIO_6 => s_writedata_from_the_iobusMDIO_6,
      s_writedata_from_the_iobusMDIO_7 => s_writedata_from_the_iobusMDIO_7,
      s_writedata_from_the_iobusREGFILE_0 => s_writedata_from_the_iobusREGFILE_0,
      txd_from_the_rs232_uart => txd_from_the_rs232_uart,
      clk1 => clk1,
      reset_n => reset_n,
      rxd_to_the_rs232_uart => rxd_to_the_rs232_uart,
      s_readdata_to_the_iobusMAC_0 => s_readdata_to_the_iobusMAC_0,
      s_readdata_to_the_iobusMAC_1 => s_readdata_to_the_iobusMAC_1,
      s_readdata_to_the_iobusMAC_2 => s_readdata_to_the_iobusMAC_2,
      s_readdata_to_the_iobusMAC_3 => s_readdata_to_the_iobusMAC_3,
      s_readdata_to_the_iobusMAC_4 => s_readdata_to_the_iobusMAC_4,
      s_readdata_to_the_iobusMAC_5 => s_readdata_to_the_iobusMAC_5,
      s_readdata_to_the_iobusMAC_6 => s_readdata_to_the_iobusMAC_6,
      s_readdata_to_the_iobusMAC_7 => s_readdata_to_the_iobusMAC_7,
      s_readdata_to_the_iobusMDIO_0 => s_readdata_to_the_iobusMDIO_0,
      s_readdata_to_the_iobusMDIO_1 => s_readdata_to_the_iobusMDIO_1,
      s_readdata_to_the_iobusMDIO_2 => s_readdata_to_the_iobusMDIO_2,
      s_readdata_to_the_iobusMDIO_3 => s_readdata_to_the_iobusMDIO_3,
      s_readdata_to_the_iobusMDIO_4 => s_readdata_to_the_iobusMDIO_4,
      s_readdata_to_the_iobusMDIO_5 => s_readdata_to_the_iobusMDIO_5,
      s_readdata_to_the_iobusMDIO_6 => s_readdata_to_the_iobusMDIO_6,
      s_readdata_to_the_iobusMDIO_7 => s_readdata_to_the_iobusMDIO_7,
      s_readdata_to_the_iobusREGFILE_0 => s_readdata_to_the_iobusREGFILE_0,
      s_readdatavalid_to_the_iobusMAC_0 => s_readdatavalid_to_the_iobusMAC_0,
      s_readdatavalid_to_the_iobusMAC_1 => s_readdatavalid_to_the_iobusMAC_1,
      s_readdatavalid_to_the_iobusMAC_2 => s_readdatavalid_to_the_iobusMAC_2,
      s_readdatavalid_to_the_iobusMAC_3 => s_readdatavalid_to_the_iobusMAC_3,
      s_readdatavalid_to_the_iobusMAC_4 => s_readdatavalid_to_the_iobusMAC_4,
      s_readdatavalid_to_the_iobusMAC_5 => s_readdatavalid_to_the_iobusMAC_5,
      s_readdatavalid_to_the_iobusMAC_6 => s_readdatavalid_to_the_iobusMAC_6,
      s_readdatavalid_to_the_iobusMAC_7 => s_readdatavalid_to_the_iobusMAC_7,
      s_readdatavalid_to_the_iobusMDIO_0 => s_readdatavalid_to_the_iobusMDIO_0,
      s_readdatavalid_to_the_iobusMDIO_1 => s_readdatavalid_to_the_iobusMDIO_1,
      s_readdatavalid_to_the_iobusMDIO_2 => s_readdatavalid_to_the_iobusMDIO_2,
      s_readdatavalid_to_the_iobusMDIO_3 => s_readdatavalid_to_the_iobusMDIO_3,
      s_readdatavalid_to_the_iobusMDIO_4 => s_readdatavalid_to_the_iobusMDIO_4,
      s_readdatavalid_to_the_iobusMDIO_5 => s_readdatavalid_to_the_iobusMDIO_5,
      s_readdatavalid_to_the_iobusMDIO_6 => s_readdatavalid_to_the_iobusMDIO_6,
      s_readdatavalid_to_the_iobusMDIO_7 => s_readdatavalid_to_the_iobusMDIO_7,
      s_readdatavalid_to_the_iobusREGFILE_0 => s_readdatavalid_to_the_iobusREGFILE_0,
      s_waitrequest_to_the_iobusMAC_0 => s_waitrequest_to_the_iobusMAC_0,
      s_waitrequest_to_the_iobusMAC_1 => s_waitrequest_to_the_iobusMAC_1,
      s_waitrequest_to_the_iobusMAC_2 => s_waitrequest_to_the_iobusMAC_2,
      s_waitrequest_to_the_iobusMAC_3 => s_waitrequest_to_the_iobusMAC_3,
      s_waitrequest_to_the_iobusMAC_4 => s_waitrequest_to_the_iobusMAC_4,
      s_waitrequest_to_the_iobusMAC_5 => s_waitrequest_to_the_iobusMAC_5,
      s_waitrequest_to_the_iobusMAC_6 => s_waitrequest_to_the_iobusMAC_6,
      s_waitrequest_to_the_iobusMAC_7 => s_waitrequest_to_the_iobusMAC_7,
      s_waitrequest_to_the_iobusMDIO_0 => s_waitrequest_to_the_iobusMDIO_0,
      s_waitrequest_to_the_iobusMDIO_1 => s_waitrequest_to_the_iobusMDIO_1,
      s_waitrequest_to_the_iobusMDIO_2 => s_waitrequest_to_the_iobusMDIO_2,
      s_waitrequest_to_the_iobusMDIO_3 => s_waitrequest_to_the_iobusMDIO_3,
      s_waitrequest_to_the_iobusMDIO_4 => s_waitrequest_to_the_iobusMDIO_4,
      s_waitrequest_to_the_iobusMDIO_5 => s_waitrequest_to_the_iobusMDIO_5,
      s_waitrequest_to_the_iobusMDIO_6 => s_waitrequest_to_the_iobusMDIO_6,
      s_waitrequest_to_the_iobusMDIO_7 => s_waitrequest_to_the_iobusMDIO_7,
      s_waitrequest_to_the_iobusREGFILE_0 => s_waitrequest_to_the_iobusREGFILE_0
    );


