// usb_control.v

// Generated using ACDS version 12.0 178 at 2012.10.18.10:39:32

`timescale 1 ps / 1 ps
module usb_control (
		output wire        m_we_from_the_ports,        // portmux.we
		output wire        m_re_from_the_ports,        //        .re
		output wire [31:0] m_writedata_from_the_ports, //        .writedata
		input  wire [31:0] m_readdata_to_the_ports,    //        .readdata
		output wire        m_reset_n_from_the_ports,   //        .reset_n
		output wire [3:0]  m_address_from_the_ports,   //        .address
		input  wire        reset_n,                    //   reset.reset_n
		output wire        CS_N_from_the_ISP1761,      //     usb.CS_N
		output wire        WR_N_from_the_ISP1761,      //        .WR_N
		output wire        RD_N_from_the_ISP1761,      //        .RD_N
		inout  wire [31:0] D_to_and_from_the_ISP1761,  //        .D
		output wire [16:0] A_from_the_ISP1761,         //        .A
		input  wire        DC_IRQ_to_the_ISP1761,      //        .DC_IRQ
		input  wire        DC_DREQ_to_the_ISP1761,     //        .DC_DREQ
		input  wire        HC_DREQ_to_the_ISP1761,     //        .HC_DREQ
		output wire        DC_DACK_from_the_ISP1761,   //        .DC_DACK
		output wire        HC_DACK_from_the_ISP1761,   //        .HC_DACK
		input  wire        HC_IRQ_to_the_ISP1761,      //        .HC_IRQ
		output wire        RESET_N_from_the_ISP1761,   //        .RESET_N
		input  wire        clk                         //     clk.clk
	);

	wire         cpu_data_master_waitrequest;                                                                 // cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                                                   // cpu:d_writedata -> cpu_data_master_translator:av_writedata
	wire  [20:0] cpu_data_master_address;                                                                     // cpu:d_address -> cpu_data_master_translator:av_address
	wire         cpu_data_master_write;                                                                       // cpu:d_write -> cpu_data_master_translator:av_write
	wire         cpu_data_master_read;                                                                        // cpu:d_read -> cpu_data_master_translator:av_read
	wire  [31:0] cpu_data_master_readdata;                                                                    // cpu_data_master_translator:av_readdata -> cpu:d_readdata
	wire   [3:0] cpu_data_master_byteenable;                                                                  // cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	wire  [31:0] isp1761_slave_translator_avalon_anti_slave_0_writedata;                                      // ISP1761_slave_translator:av_writedata -> ISP1761:s_writedata
	wire  [17:0] isp1761_slave_translator_avalon_anti_slave_0_address;                                        // ISP1761_slave_translator:av_address -> ISP1761:s_address
	wire         isp1761_slave_translator_avalon_anti_slave_0_chipselect;                                     // ISP1761_slave_translator:av_chipselect -> ISP1761:s_cs_n
	wire         isp1761_slave_translator_avalon_anti_slave_0_write;                                          // ISP1761_slave_translator:av_write -> ISP1761:s_write_n
	wire         isp1761_slave_translator_avalon_anti_slave_0_read;                                           // ISP1761_slave_translator:av_read -> ISP1761:s_read_n
	wire  [31:0] isp1761_slave_translator_avalon_anti_slave_0_readdata;                                       // ISP1761:s_readdata -> ISP1761_slave_translator:av_readdata
	wire  [31:0] ports_slave_translator_avalon_anti_slave_0_writedata;                                        // ports_slave_translator:av_writedata -> ports:s_writedata
	wire   [3:0] ports_slave_translator_avalon_anti_slave_0_address;                                          // ports_slave_translator:av_address -> ports:s_address
	wire         ports_slave_translator_avalon_anti_slave_0_write;                                            // ports_slave_translator:av_write -> ports:s_we
	wire         ports_slave_translator_avalon_anti_slave_0_read;                                             // ports_slave_translator:av_read -> ports:s_re
	wire  [31:0] ports_slave_translator_avalon_anti_slave_0_readdata;                                         // ports:s_readdata -> ports_slave_translator:av_readdata
	wire         cpu_tightly_coupled_instruction_master_0_waitrequest;                                        // cpu_tightly_coupled_instruction_master_0_translator:av_waitrequest -> cpu:icm0_waitrequest
	wire  [22:0] cpu_tightly_coupled_instruction_master_0_address;                                            // cpu:icm0_address -> cpu_tightly_coupled_instruction_master_0_translator:av_address
	wire         cpu_tightly_coupled_instruction_master_0_clken;                                              // cpu:icm0_clken -> cpu_tightly_coupled_instruction_master_0_translator:av_clken
	wire         cpu_tightly_coupled_instruction_master_0_read;                                               // cpu:icm0_read -> cpu_tightly_coupled_instruction_master_0_translator:av_read
	wire  [31:0] cpu_tightly_coupled_instruction_master_0_readdata;                                           // cpu_tightly_coupled_instruction_master_0_translator:av_readdata -> cpu:icm0_readdata
	wire         cpu_tightly_coupled_instruction_master_0_readdatavalid;                                      // cpu_tightly_coupled_instruction_master_0_translator:av_readdatavalid -> cpu:icm0_readdatavalid
	wire         cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_waitrequest;   // mem_s1_translator:uav_waitrequest -> cpu_tightly_coupled_instruction_master_0_translator:uav_waitrequest
	wire   [2:0] cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_burstcount;    // cpu_tightly_coupled_instruction_master_0_translator:uav_burstcount -> mem_s1_translator:uav_burstcount
	wire  [31:0] cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_writedata;     // cpu_tightly_coupled_instruction_master_0_translator:uav_writedata -> mem_s1_translator:uav_writedata
	wire  [22:0] cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_address;       // cpu_tightly_coupled_instruction_master_0_translator:uav_address -> mem_s1_translator:uav_address
	wire         cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_clken;         // cpu_tightly_coupled_instruction_master_0_translator:uav_clken -> mem_s1_translator:uav_clken
	wire         cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_lock;          // cpu_tightly_coupled_instruction_master_0_translator:uav_lock -> mem_s1_translator:uav_lock
	wire         cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_write;         // cpu_tightly_coupled_instruction_master_0_translator:uav_write -> mem_s1_translator:uav_write
	wire         cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_read;          // cpu_tightly_coupled_instruction_master_0_translator:uav_read -> mem_s1_translator:uav_read
	wire  [31:0] cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_readdata;      // mem_s1_translator:uav_readdata -> cpu_tightly_coupled_instruction_master_0_translator:uav_readdata
	wire         cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_debugaccess;   // cpu_tightly_coupled_instruction_master_0_translator:uav_debugaccess -> mem_s1_translator:uav_debugaccess
	wire   [3:0] cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_byteenable;    // cpu_tightly_coupled_instruction_master_0_translator:uav_byteenable -> mem_s1_translator:uav_byteenable
	wire         cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_readdatavalid; // mem_s1_translator:uav_readdatavalid -> cpu_tightly_coupled_instruction_master_0_translator:uav_readdatavalid
	wire  [31:0] mem_s1_translator_avalon_anti_slave_0_writedata;                                             // mem_s1_translator:av_writedata -> mem:writedata
	wire  [10:0] mem_s1_translator_avalon_anti_slave_0_address;                                               // mem_s1_translator:av_address -> mem:address
	wire         mem_s1_translator_avalon_anti_slave_0_chipselect;                                            // mem_s1_translator:av_chipselect -> mem:chipselect
	wire         mem_s1_translator_avalon_anti_slave_0_clken;                                                 // mem_s1_translator:av_clken -> mem:clken
	wire         mem_s1_translator_avalon_anti_slave_0_write;                                                 // mem_s1_translator:av_write -> mem:write
	wire  [31:0] mem_s1_translator_avalon_anti_slave_0_readdata;                                              // mem:readdata -> mem_s1_translator:av_readdata
	wire   [3:0] mem_s1_translator_avalon_anti_slave_0_byteenable;                                            // mem_s1_translator:av_byteenable -> mem:byteenable
	wire         cpu_tightly_coupled_data_master_0_waitrequest;                                               // cpu_tightly_coupled_data_master_0_translator:av_waitrequest -> cpu:dcm0_waitrequest
	wire  [31:0] cpu_tightly_coupled_data_master_0_writedata;                                                 // cpu:dcm0_writedata -> cpu_tightly_coupled_data_master_0_translator:av_writedata
	wire  [22:0] cpu_tightly_coupled_data_master_0_address;                                                   // cpu:dcm0_address -> cpu_tightly_coupled_data_master_0_translator:av_address
	wire         cpu_tightly_coupled_data_master_0_clken;                                                     // cpu:dcm0_clken -> cpu_tightly_coupled_data_master_0_translator:av_clken
	wire         cpu_tightly_coupled_data_master_0_write;                                                     // cpu:dcm0_write -> cpu_tightly_coupled_data_master_0_translator:av_write
	wire         cpu_tightly_coupled_data_master_0_read;                                                      // cpu:dcm0_read -> cpu_tightly_coupled_data_master_0_translator:av_read
	wire  [31:0] cpu_tightly_coupled_data_master_0_readdata;                                                  // cpu_tightly_coupled_data_master_0_translator:av_readdata -> cpu:dcm0_readdata
	wire   [3:0] cpu_tightly_coupled_data_master_0_byteenable;                                                // cpu:dcm0_byteenable -> cpu_tightly_coupled_data_master_0_translator:av_byteenable
	wire         cpu_tightly_coupled_data_master_0_readdatavalid;                                             // cpu_tightly_coupled_data_master_0_translator:av_readdatavalid -> cpu:dcm0_readdatavalid
	wire         cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_waitrequest;          // mem_s2_translator:uav_waitrequest -> cpu_tightly_coupled_data_master_0_translator:uav_waitrequest
	wire   [2:0] cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_burstcount;           // cpu_tightly_coupled_data_master_0_translator:uav_burstcount -> mem_s2_translator:uav_burstcount
	wire  [31:0] cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_writedata;            // cpu_tightly_coupled_data_master_0_translator:uav_writedata -> mem_s2_translator:uav_writedata
	wire  [22:0] cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_address;              // cpu_tightly_coupled_data_master_0_translator:uav_address -> mem_s2_translator:uav_address
	wire         cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_clken;                // cpu_tightly_coupled_data_master_0_translator:uav_clken -> mem_s2_translator:uav_clken
	wire         cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_lock;                 // cpu_tightly_coupled_data_master_0_translator:uav_lock -> mem_s2_translator:uav_lock
	wire         cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_write;                // cpu_tightly_coupled_data_master_0_translator:uav_write -> mem_s2_translator:uav_write
	wire         cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_read;                 // cpu_tightly_coupled_data_master_0_translator:uav_read -> mem_s2_translator:uav_read
	wire  [31:0] cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_readdata;             // mem_s2_translator:uav_readdata -> cpu_tightly_coupled_data_master_0_translator:uav_readdata
	wire         cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_debugaccess;          // cpu_tightly_coupled_data_master_0_translator:uav_debugaccess -> mem_s2_translator:uav_debugaccess
	wire   [3:0] cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_byteenable;           // cpu_tightly_coupled_data_master_0_translator:uav_byteenable -> mem_s2_translator:uav_byteenable
	wire         cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_readdatavalid;        // mem_s2_translator:uav_readdatavalid -> cpu_tightly_coupled_data_master_0_translator:uav_readdatavalid
	wire  [31:0] mem_s2_translator_avalon_anti_slave_0_writedata;                                             // mem_s2_translator:av_writedata -> mem:writedata2
	wire  [10:0] mem_s2_translator_avalon_anti_slave_0_address;                                               // mem_s2_translator:av_address -> mem:address2
	wire         mem_s2_translator_avalon_anti_slave_0_chipselect;                                            // mem_s2_translator:av_chipselect -> mem:chipselect2
	wire         mem_s2_translator_avalon_anti_slave_0_clken;                                                 // mem_s2_translator:av_clken -> mem:clken2
	wire         mem_s2_translator_avalon_anti_slave_0_write;                                                 // mem_s2_translator:av_write -> mem:write2
	wire  [31:0] mem_s2_translator_avalon_anti_slave_0_readdata;                                              // mem:readdata2 -> mem_s2_translator:av_readdata
	wire   [3:0] mem_s2_translator_avalon_anti_slave_0_byteenable;                                            // mem_s2_translator:av_byteenable -> mem:byteenable2
	wire         cpu_data_master_translator_avalon_universal_master_0_waitrequest;                            // cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	wire   [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                             // cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                              // cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [20:0] cpu_data_master_translator_avalon_universal_master_0_address;                                // cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         cpu_data_master_translator_avalon_universal_master_0_lock;                                   // cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         cpu_data_master_translator_avalon_universal_master_0_write;                                  // cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         cpu_data_master_translator_avalon_universal_master_0_read;                                   // cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                               // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	wire         cpu_data_master_translator_avalon_universal_master_0_debugaccess;                            // cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                             // cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                          // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // ISP1761_slave_translator:uav_waitrequest -> ISP1761_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] isp1761_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // ISP1761_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> ISP1761_slave_translator:uav_burstcount
	wire  [31:0] isp1761_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                        // ISP1761_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> ISP1761_slave_translator:uav_writedata
	wire  [20:0] isp1761_slave_translator_avalon_universal_slave_0_agent_m0_address;                          // ISP1761_slave_translator_avalon_universal_slave_0_agent:m0_address -> ISP1761_slave_translator:uav_address
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_m0_write;                            // ISP1761_slave_translator_avalon_universal_slave_0_agent:m0_write -> ISP1761_slave_translator:uav_write
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_m0_lock;                             // ISP1761_slave_translator_avalon_universal_slave_0_agent:m0_lock -> ISP1761_slave_translator:uav_lock
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_m0_read;                             // ISP1761_slave_translator_avalon_universal_slave_0_agent:m0_read -> ISP1761_slave_translator:uav_read
	wire  [31:0] isp1761_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                         // ISP1761_slave_translator:uav_readdata -> ISP1761_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // ISP1761_slave_translator:uav_readdatavalid -> ISP1761_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // ISP1761_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ISP1761_slave_translator:uav_debugaccess
	wire   [3:0] isp1761_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // ISP1761_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> ISP1761_slave_translator:uav_byteenable
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // ISP1761_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ISP1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // ISP1761_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> ISP1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // ISP1761_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ISP1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [88:0] isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                      // ISP1761_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> ISP1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // ISP1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ISP1761_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // ISP1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ISP1761_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // ISP1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ISP1761_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // ISP1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ISP1761_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [88:0] isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // ISP1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ISP1761_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // ISP1761_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ISP1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // ISP1761_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ISP1761_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] isp1761_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // ISP1761_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ISP1761_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // ISP1761_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ISP1761_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         ports_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // ports_slave_translator:uav_waitrequest -> ports_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] ports_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // ports_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> ports_slave_translator:uav_burstcount
	wire  [31:0] ports_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // ports_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> ports_slave_translator:uav_writedata
	wire  [20:0] ports_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // ports_slave_translator_avalon_universal_slave_0_agent:m0_address -> ports_slave_translator:uav_address
	wire         ports_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // ports_slave_translator_avalon_universal_slave_0_agent:m0_write -> ports_slave_translator:uav_write
	wire         ports_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // ports_slave_translator_avalon_universal_slave_0_agent:m0_lock -> ports_slave_translator:uav_lock
	wire         ports_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // ports_slave_translator_avalon_universal_slave_0_agent:m0_read -> ports_slave_translator:uav_read
	wire  [31:0] ports_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // ports_slave_translator:uav_readdata -> ports_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         ports_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // ports_slave_translator:uav_readdatavalid -> ports_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         ports_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // ports_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ports_slave_translator:uav_debugaccess
	wire   [3:0] ports_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // ports_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> ports_slave_translator:uav_byteenable
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // ports_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // ports_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // ports_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [88:0] ports_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // ports_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ports_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ports_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ports_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ports_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [88:0] ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ports_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // ports_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // ports_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ports_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] ports_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // ports_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ports_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // ports_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ports_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                   // cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                         // cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                 // cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [87:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                          // cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                         // addr_router:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // ISP1761_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rp_valid;                            // ISP1761_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // ISP1761_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [87:0] isp1761_slave_translator_avalon_universal_slave_0_agent_rp_data;                             // ISP1761_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         isp1761_slave_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router:sink_ready -> ISP1761_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // ports_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // ports_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // ports_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [87:0] ports_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // ports_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         ports_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_001:sink_ready -> ports_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         rst_controller_reset_out_reset;                                                              // rst_controller:reset_out -> [ISP1761:s_reset_n, ISP1761_slave_translator:reset, ISP1761_slave_translator_avalon_universal_slave_0_agent:reset, ISP1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, cmd_xbar_demux:reset, cpu:reset_n, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_tightly_coupled_data_master_0_translator:reset, cpu_tightly_coupled_instruction_master_0_translator:reset, id_router:reset, id_router_001:reset, irq_mapper:reset, mem:reset, mem:reset2, mem_s1_translator:reset, mem_s2_translator:reset, ports:s_reset_n, ports_slave_translator:reset, ports_slave_translator_avalon_universal_slave_0_agent:reset, ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_mux:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                             // cmd_xbar_demux:src0_endofpacket -> ISP1761_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                   // cmd_xbar_demux:src0_valid -> ISP1761_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                           // cmd_xbar_demux:src0_startofpacket -> ISP1761_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [87:0] cmd_xbar_demux_src0_data;                                                                    // cmd_xbar_demux:src0_data -> ISP1761_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_demux_src0_channel;                                                                 // cmd_xbar_demux:src0_channel -> ISP1761_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_src1_endofpacket;                                                             // cmd_xbar_demux:src1_endofpacket -> ports_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                   // cmd_xbar_demux:src1_valid -> ports_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                           // cmd_xbar_demux:src1_startofpacket -> ports_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [87:0] cmd_xbar_demux_src1_data;                                                                    // cmd_xbar_demux:src1_data -> ports_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [1:0] cmd_xbar_demux_src1_channel;                                                                 // cmd_xbar_demux:src1_channel -> ports_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                             // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                   // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                           // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [87:0] rsp_xbar_demux_src0_data;                                                                    // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [1:0] rsp_xbar_demux_src0_channel;                                                                 // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                   // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                         // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                               // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                       // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [87:0] rsp_xbar_demux_001_src0_data;                                                                // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire   [1:0] rsp_xbar_demux_001_src0_channel;                                                             // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                               // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         addr_router_src_endofpacket;                                                                 // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         addr_router_src_valid;                                                                       // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire         addr_router_src_startofpacket;                                                               // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [87:0] addr_router_src_data;                                                                        // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [1:0] addr_router_src_channel;                                                                     // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire         addr_router_src_ready;                                                                       // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                // rsp_xbar_mux:src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                      // rsp_xbar_mux:src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                              // rsp_xbar_mux:src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [87:0] rsp_xbar_mux_src_data;                                                                       // rsp_xbar_mux:src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [1:0] rsp_xbar_mux_src_channel;                                                                    // rsp_xbar_mux:src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         rsp_xbar_mux_src_ready;                                                                      // cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire         cmd_xbar_demux_src0_ready;                                                                   // ISP1761_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src0_ready
	wire         id_router_src_endofpacket;                                                                   // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                         // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                 // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [87:0] id_router_src_data;                                                                          // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [1:0] id_router_src_channel;                                                                       // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                         // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_demux_src1_ready;                                                                   // ports_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src1_ready
	wire         id_router_001_src_endofpacket;                                                               // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                     // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                             // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [87:0] id_router_001_src_data;                                                                      // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [1:0] id_router_001_src_channel;                                                                   // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                     // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire  [31:0] cpu_d_irq_irq;                                                                               // irq_mapper:sender_irq -> cpu:d_irq

	usb_control_mem mem (
		.clk         (clk),                                              //   clk1.clk
		.address     (mem_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect  (mem_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken       (mem_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata    (mem_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write       (mem_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata   (mem_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable  (mem_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                   // reset1.reset
		.address2    (mem_s2_translator_avalon_anti_slave_0_address),    //     s2.address
		.chipselect2 (mem_s2_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken2      (mem_s2_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata2   (mem_s2_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write2      (mem_s2_translator_avalon_anti_slave_0_write),      //       .write
		.writedata2  (mem_s2_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable2 (mem_s2_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.clk2        (clk),                                              //   clk2.clk
		.reset2      (rst_controller_reset_out_reset)                    // reset2.reset
	);

	ISP1761_IF isp1761 (
		.CS_N        (CS_N_from_the_ISP1761),                                    //       usb.export
		.WR_N        (WR_N_from_the_ISP1761),                                    //          .export
		.RD_N        (RD_N_from_the_ISP1761),                                    //          .export
		.D           (D_to_and_from_the_ISP1761),                                //          .export
		.A           (A_from_the_ISP1761),                                       //          .export
		.DC_IRQ      (DC_IRQ_to_the_ISP1761),                                    //          .export
		.DC_DREQ     (DC_DREQ_to_the_ISP1761),                                   //          .export
		.HC_DREQ     (HC_DREQ_to_the_ISP1761),                                   //          .export
		.DC_DACK     (DC_DACK_from_the_ISP1761),                                 //          .export
		.HC_DACK     (HC_DACK_from_the_ISP1761),                                 //          .export
		.HC_IRQ      (HC_IRQ_to_the_ISP1761),                                    //          .export
		.RESET_N     (RESET_N_from_the_ISP1761),                                 //          .export
		.s_address   (isp1761_slave_translator_avalon_anti_slave_0_address),     //     slave.address
		.s_write_n   (~isp1761_slave_translator_avalon_anti_slave_0_write),      //          .write_n
		.s_writedata (isp1761_slave_translator_avalon_anti_slave_0_writedata),   //          .writedata
		.s_read_n    (~isp1761_slave_translator_avalon_anti_slave_0_read),       //          .read_n
		.s_readdata  (isp1761_slave_translator_avalon_anti_slave_0_readdata),    //          .readdata
		.s_cs_n      (~isp1761_slave_translator_avalon_anti_slave_0_chipselect), //          .chipselect_n
		.s_irq       (),                                                         // slave_irq.irq
		.s_clk       (clk),                                                      //       clk.clk
		.s_reset_n   (~rst_controller_reset_out_reset)                           //     reset.reset_n
	);

	portmux_export ports (
		.s_we        (ports_slave_translator_avalon_anti_slave_0_write),     //  slave.write
		.s_re        (ports_slave_translator_avalon_anti_slave_0_read),      //       .read
		.s_writedata (ports_slave_translator_avalon_anti_slave_0_writedata), //       .writedata
		.s_readdata  (ports_slave_translator_avalon_anti_slave_0_readdata),  //       .readdata
		.s_address   (ports_slave_translator_avalon_anti_slave_0_address),   //       .address
		.m_we        (m_we_from_the_ports),                                  // export.export
		.m_re        (m_re_from_the_ports),                                  //       .export
		.m_writedata (m_writedata_from_the_ports),                           //       .export
		.m_readdata  (m_readdata_to_the_ports),                              //       .export
		.m_reset_n   (m_reset_n_from_the_ports),                             //       .export
		.m_address   (m_address_from_the_ports),                             //       .export
		.s_reset_n   (~rst_controller_reset_out_reset),                      //  reset.reset_n
		.s_clk       (clk)                                                   //    clk.clk
	);

	usb_control_cpu cpu (
		.clk                (clk),                                                    //                                  clk.clk
		.reset_n            (~rst_controller_reset_out_reset),                        //                              reset_n.reset_n
		.d_address          (cpu_data_master_address),                                //                          data_master.address
		.d_byteenable       (cpu_data_master_byteenable),                             //                                     .byteenable
		.d_read             (cpu_data_master_read),                                   //                                     .read
		.d_readdata         (cpu_data_master_readdata),                               //                                     .readdata
		.d_waitrequest      (cpu_data_master_waitrequest),                            //                                     .waitrequest
		.d_write            (cpu_data_master_write),                                  //                                     .write
		.d_writedata        (cpu_data_master_writedata),                              //                                     .writedata
		.dcm0_readdata      (cpu_tightly_coupled_data_master_0_readdata),             //        tightly_coupled_data_master_0.readdata
		.dcm0_waitrequest   (cpu_tightly_coupled_data_master_0_waitrequest),          //                                     .waitrequest
		.dcm0_readdatavalid (cpu_tightly_coupled_data_master_0_readdatavalid),        //                                     .readdatavalid
		.dcm0_address       (cpu_tightly_coupled_data_master_0_address),              //                                     .address
		.dcm0_read          (cpu_tightly_coupled_data_master_0_read),                 //                                     .read
		.dcm0_clken         (cpu_tightly_coupled_data_master_0_clken),                //                                     .clken
		.dcm0_byteenable    (cpu_tightly_coupled_data_master_0_byteenable),           //                                     .byteenable
		.dcm0_write         (cpu_tightly_coupled_data_master_0_write),                //                                     .write
		.dcm0_writedata     (cpu_tightly_coupled_data_master_0_writedata),            //                                     .writedata
		.icm0_readdata      (cpu_tightly_coupled_instruction_master_0_readdata),      // tightly_coupled_instruction_master_0.readdata
		.icm0_waitrequest   (cpu_tightly_coupled_instruction_master_0_waitrequest),   //                                     .waitrequest
		.icm0_readdatavalid (cpu_tightly_coupled_instruction_master_0_readdatavalid), //                                     .readdatavalid
		.icm0_address       (cpu_tightly_coupled_instruction_master_0_address),       //                                     .address
		.icm0_read          (cpu_tightly_coupled_instruction_master_0_read),          //                                     .read
		.icm0_clken         (cpu_tightly_coupled_instruction_master_0_clken),         //                                     .clken
		.d_irq              (cpu_d_irq_irq),                                          //                                d_irq.irq
		.no_ci_readra       ()                                                        //            custom_instruction_master.readra
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (21),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (21),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_data_master_translator (
		.clk                   (clk),                                                                //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address           (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read               (cpu_data_master_read),                                               //                          .read
		.av_readdata           (cpu_data_master_readdata),                                           //                          .readdata
		.av_write              (cpu_data_master_write),                                              //                          .write
		.av_writedata          (cpu_data_master_writedata),                                          //                          .writedata
		.av_burstcount         (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer (1'b0),                                                               //               (terminated)
		.av_begintransfer      (1'b0),                                                               //               (terminated)
		.av_chipselect         (1'b0),                                                               //               (terminated)
		.av_readdatavalid      (),                                                                   //               (terminated)
		.av_lock               (1'b0),                                                               //               (terminated)
		.av_debugaccess        (1'b0),                                                               //               (terminated)
		.uav_clken             (),                                                                   //               (terminated)
		.av_clken              (1'b1)                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (18),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (2),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (1),
		.AV_DATA_HOLD_CYCLES            (1)
	) isp1761_slave_translator (
		.clk                   (clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (isp1761_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (isp1761_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (isp1761_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (isp1761_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (isp1761_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (isp1761_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (4),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ports_slave_translator (
		.clk                   (clk),                                                                    //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address           (ports_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (ports_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (ports_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (ports_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (ports_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (ports_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (ports_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (ports_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (ports_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (ports_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (ports_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (ports_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (ports_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (ports_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (ports_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (ports_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_chipselect         (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (23),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (23),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_tightly_coupled_instruction_master_0_translator (
		.clk                   (clk),                                                                                         //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                              //                     reset.reset
		.uav_address           (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.uav_clken             (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_clken),         //                          .clken
		.av_address            (cpu_tightly_coupled_instruction_master_0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_tightly_coupled_instruction_master_0_waitrequest),                                        //                          .waitrequest
		.av_read               (cpu_tightly_coupled_instruction_master_0_read),                                               //                          .read
		.av_readdata           (cpu_tightly_coupled_instruction_master_0_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_tightly_coupled_instruction_master_0_readdatavalid),                                      //                          .readdatavalid
		.av_clken              (cpu_tightly_coupled_instruction_master_0_clken),                                              //                          .clken
		.av_burstcount         (1'b1),                                                                                        //               (terminated)
		.av_byteenable         (4'b1111),                                                                                     //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                        //               (terminated)
		.av_begintransfer      (1'b0),                                                                                        //               (terminated)
		.av_chipselect         (1'b0),                                                                                        //               (terminated)
		.av_write              (1'b0),                                                                                        //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                                        //               (terminated)
		.av_lock               (1'b0),                                                                                        //               (terminated)
		.av_debugaccess        (1'b0)                                                                                         //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (23),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (1),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mem_s1_translator (
		.clk                   (clk),                                                                                         //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                              //                    reset.reset
		.uav_address           (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read              (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write             (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest       (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata         (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock              (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess       (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.uav_clken             (cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_clken),         //                         .clken
		.av_address            (mem_s1_translator_avalon_anti_slave_0_address),                                               //      avalon_anti_slave_0.address
		.av_write              (mem_s1_translator_avalon_anti_slave_0_write),                                                 //                         .write
		.av_readdata           (mem_s1_translator_avalon_anti_slave_0_readdata),                                              //                         .readdata
		.av_writedata          (mem_s1_translator_avalon_anti_slave_0_writedata),                                             //                         .writedata
		.av_byteenable         (mem_s1_translator_avalon_anti_slave_0_byteenable),                                            //                         .byteenable
		.av_chipselect         (mem_s1_translator_avalon_anti_slave_0_chipselect),                                            //                         .chipselect
		.av_clken              (mem_s1_translator_avalon_anti_slave_0_clken),                                                 //                         .clken
		.av_read               (),                                                                                            //              (terminated)
		.av_begintransfer      (),                                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                                            //              (terminated)
		.av_burstcount         (),                                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                                            //              (terminated)
		.av_lock               (),                                                                                            //              (terminated)
		.av_debugaccess        (),                                                                                            //              (terminated)
		.av_outputenable       ()                                                                                             //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (23),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (23),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_tightly_coupled_data_master_0_translator (
		.clk                   (clk),                                                                                  //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                       //                     reset.reset
		.uav_address           (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.uav_clken             (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_clken),         //                          .clken
		.av_address            (cpu_tightly_coupled_data_master_0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (cpu_tightly_coupled_data_master_0_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (cpu_tightly_coupled_data_master_0_byteenable),                                         //                          .byteenable
		.av_read               (cpu_tightly_coupled_data_master_0_read),                                               //                          .read
		.av_readdata           (cpu_tightly_coupled_data_master_0_readdata),                                           //                          .readdata
		.av_readdatavalid      (cpu_tightly_coupled_data_master_0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (cpu_tightly_coupled_data_master_0_write),                                              //                          .write
		.av_writedata          (cpu_tightly_coupled_data_master_0_writedata),                                          //                          .writedata
		.av_clken              (cpu_tightly_coupled_data_master_0_clken),                                              //                          .clken
		.av_burstcount         (1'b1),                                                                                 //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                                 //               (terminated)
		.av_begintransfer      (1'b0),                                                                                 //               (terminated)
		.av_chipselect         (1'b0),                                                                                 //               (terminated)
		.av_lock               (1'b0),                                                                                 //               (terminated)
		.av_debugaccess        (1'b0)                                                                                  //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (23),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (1),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) mem_s2_translator (
		.clk                   (clk),                                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                       //                    reset.reset
		.uav_address           (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_burstcount),    //                         .burstcount
		.uav_read              (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_read),          //                         .read
		.uav_write             (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_write),         //                         .write
		.uav_waitrequest       (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_byteenable),    //                         .byteenable
		.uav_readdata          (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_readdata),      //                         .readdata
		.uav_writedata         (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_writedata),     //                         .writedata
		.uav_lock              (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_lock),          //                         .lock
		.uav_debugaccess       (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_debugaccess),   //                         .debugaccess
		.uav_clken             (cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_clken),         //                         .clken
		.av_address            (mem_s2_translator_avalon_anti_slave_0_address),                                        //      avalon_anti_slave_0.address
		.av_write              (mem_s2_translator_avalon_anti_slave_0_write),                                          //                         .write
		.av_readdata           (mem_s2_translator_avalon_anti_slave_0_readdata),                                       //                         .readdata
		.av_writedata          (mem_s2_translator_avalon_anti_slave_0_writedata),                                      //                         .writedata
		.av_byteenable         (mem_s2_translator_avalon_anti_slave_0_byteenable),                                     //                         .byteenable
		.av_chipselect         (mem_s2_translator_avalon_anti_slave_0_chipselect),                                     //                         .chipselect
		.av_clken              (mem_s2_translator_avalon_anti_slave_0_clken),                                          //                         .clken
		.av_read               (),                                                                                     //              (terminated)
		.av_begintransfer      (),                                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                                     //              (terminated)
		.av_burstcount         (),                                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                                     //              (terminated)
		.av_lock               (),                                                                                     //              (terminated)
		.av_debugaccess        (),                                                                                     //              (terminated)
		.av_outputenable       ()                                                                                      //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (79),
		.PKT_BEGIN_BURST           (75),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.PKT_BURST_TYPE_H          (73),
		.PKT_BURST_TYPE_L          (72),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_TRANS_EXCLUSIVE       (62),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (77),
		.PKT_DEST_ID_L             (77),
		.PKT_THREAD_ID_H           (78),
		.PKT_THREAD_ID_L           (78),
		.PKT_CACHE_H               (85),
		.PKT_CACHE_L               (82),
		.PKT_ADDR_SIDEBAND_H       (74),
		.PKT_ADDR_SIDEBAND_L       (74),
		.ST_DATA_W                 (88),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (4'b0000)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk),                                                                         //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address       (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (rsp_xbar_mux_src_valid),                                                      //        rp.valid
		.rp_data          (rsp_xbar_mux_src_data),                                                       //          .data
		.rp_channel       (rsp_xbar_mux_src_channel),                                                    //          .channel
		.rp_startofpacket (rsp_xbar_mux_src_startofpacket),                                              //          .startofpacket
		.rp_endofpacket   (rsp_xbar_mux_src_endofpacket),                                                //          .endofpacket
		.rp_ready         (rsp_xbar_mux_src_ready)                                                       //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (77),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (79),
		.PKT_RESPONSE_STATUS_H     (87),
		.PKT_RESPONSE_STATUS_L     (86),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (88),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) isp1761_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (isp1761_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (isp1761_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (isp1761_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (isp1761_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (isp1761_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (isp1761_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src0_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_src0_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_src0_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_src0_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src0_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src0_channel),                                                        //                .channel
		.rf_sink_ready           (isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (isp1761_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (isp1761_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (isp1761_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (isp1761_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (isp1761_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (isp1761_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (89),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (isp1761_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (isp1761_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (75),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (76),
		.PKT_SRC_ID_L              (76),
		.PKT_DEST_ID_H             (77),
		.PKT_DEST_ID_L             (77),
		.PKT_BURSTWRAP_H           (68),
		.PKT_BURSTWRAP_L           (66),
		.PKT_BYTE_CNT_H            (65),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (81),
		.PKT_PROTECTION_L          (79),
		.PKT_RESPONSE_STATUS_H     (87),
		.PKT_RESPONSE_STATUS_L     (86),
		.PKT_BURST_SIZE_H          (71),
		.PKT_BURST_SIZE_L          (69),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (88),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) ports_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (ports_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ports_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ports_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ports_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ports_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ports_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ports_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ports_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ports_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ports_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ports_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ports_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ports_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ports_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ports_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ports_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src1_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_src1_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_src1_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_src1_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src1_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src1_channel),                                                      //                .channel
		.rf_sink_ready           (ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ports_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ports_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ports_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ports_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ports_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ports_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ports_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ports_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ports_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ports_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ports_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (89),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (ports_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ports_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ports_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ports_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ports_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ports_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	usb_control_addr_router addr_router (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                       //          .valid
		.src_data           (addr_router_src_data),                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                  //          .endofpacket
	);

	usb_control_id_router id_router (
		.sink_ready         (isp1761_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (isp1761_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (isp1761_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (isp1761_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (isp1761_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                      //       src.ready
		.src_valid          (id_router_src_valid),                                                      //          .valid
		.src_data           (id_router_src_data),                                                       //          .data
		.src_channel        (id_router_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                 //          .endofpacket
	);

	usb_control_id_router id_router_001 (
		.sink_ready         (ports_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ports_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ports_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ports_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ports_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                //       src.ready
		.src_valid          (id_router_001_src_valid),                                                //          .valid
		.src_data           (id_router_001_src_data),                                                 //          .data
		.src_channel        (id_router_001_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                           //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_n),                       // reset_in0.reset
		.clk        (clk),                            //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	usb_control_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	usb_control_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)    //          .endofpacket
	);

	usb_control_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	usb_control_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk),                                   //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	usb_control_irq_mapper irq_mapper (
		.clk        (clk),                            //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (cpu_d_irq_irq)                   //    sender.irq
	);

endmodule
